//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�www.openedv.com
//�Ա����̣�http://openedv.taobao.com 
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2018-2028
//All rights reserved
//----------------------------------------------------------------------------------------
// File name:           asyn_rst_syn
// Last modified Date:  2019/7/1 9:30:00
// Last Version:        V1.1
// Descriptions:        �첽��λ��ͬ���ͷţ���ת���ɸߵ�ƽ��Ч
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2019/7/1 9:30:00
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module asyn_rst_syn(
    input clk,          //Ŀ��ʱ����
    input reset_n,      //�첽��λ������Ч
    
    output syn_reset    //����Ч
    );
    
    //reg define
    reg reset_1;
    reg reset_2;
        
    //*****************************************************
    //**                    main code
    //***************************************************** 
    assign syn_reset  = reset_2;
        
    //���첽��λ�źŽ���ͬ���ͷţ���ת���ɸ���Ч
    always @ (posedge clk or negedge reset_n) begin
        if(!reset_n) begin
            reset_1 <= 1'b1;
            reset_2 <= 1'b1;
        end
        else begin
            reset_1 <= 1'b0;
            reset_2 <= reset_1;
        end
    end
    
endmodule
